

module test();

endmodule
